// =============================================================================
// @File         :  top_test.v
// @Author       :  Jiangxuan Li
// @Created      :  2022/3/20 21:36:01
// @Description  :  top test file for modules
// 
// -----------------------------------------------------------------------------
// History
// -----------------------------------------------------------------------------
// Ver  :| Author  :| Mod. Date          :| Changes Made :|
// 0.1   | Jx L     | 2022/3/20 21:36:01 | original
// =============================================================================

module top_test (
	 input clk    // Clock
	,input rst_n
);



endmodule