// =============================================================================
// @File         :  wb_stage.v
// @Author       :  Jiangxuan Li
// @Created      :  2022/5/1 22:28:59
// @Description  :  write back stage
// 
// -----------------------------------------------------------------------------
// History
// -----------------------------------------------------------------------------
// Ver  :| Author  :| Mod. Date          :| Changes Made :|
// 0.1   | Jx L     | 2022/5/1 22:28:59 | original
// =============================================================================

module wb_stage (
	 input clk    // Clock
	,input rst_n  // Asynchronous reset active low
	,
);



endmodule
